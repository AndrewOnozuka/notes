//`include "fulladder.sv"
module carry_lookahead_adder#(parameter N=4)(
  input logic[N-1:0] A, B,
  input logic CIN,
  output logic[N:0] result
);

 // Add code for carry lookahead adder 
  
endmodule: carry_lookahead_adder

